-- defender_common: Package containing common constants for FPGA defender
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package defender_common is

    
    
    
end package defender_common;